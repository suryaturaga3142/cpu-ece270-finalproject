// Combined all ALU related things into this