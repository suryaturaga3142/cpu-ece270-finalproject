`default_nettype none
`include "params.svh"

`ifndef sequencer_guard
`define sequencer_guard

// Code here

`endif