module RAM_wrapper(

    input logic en, 
    input logic 

)



endmodule