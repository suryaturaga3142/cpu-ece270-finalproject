// Combined all ALU related things into this
`default_nettype none
`include "params.svh"
`ifndef alu_guard
`define alu_guard

module alu (
    input logic clk, rstn
    
);
    
endmodule
`endif 