module ROM(

); 



endmodule