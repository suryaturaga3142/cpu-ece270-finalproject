`include "cpu.sv"